module hexdriver (input [25:0] val, output reg [6:0] HEX1, output reg [6:0] HEX2);


	always_comb
		case(val)
		
		// Ridiculously long case statement to output proper display values
		
		// 01 ~
		26'b00000000000000000000000001: begin
		HEX1 <= 7'b100_0000; // 0
		HEX2 <= 7'b111_1001; // 1
		end
		
		// 02 ~
		26'b00000000000000000000000010: begin
		HEX1 <= 7'b100_0000; // 0
		HEX2 <= 7'b010_0100; // 2
		end
		
		// 03 ~
		26'b00000000000000000000000100: begin
		HEX1 <= 7'b100_0000; // 0
		HEX2 <= 7'b011_0000; // 3
		end
		
		// 04 ~
		26'b00000000000000000000001000: begin
		HEX1 <= 7'b100_0000;  
		HEX2 <= 7'b001_1001;
		end
		
		// 05 ~
		26'b00000000000000000000010000: begin
		HEX1 <= 7'b100_0000; // 0
		HEX2 <= 7'b001_0010; // 5
		end
		
		// 06 ~
		26'b00000000000000000000100000: begin
		HEX1 <= 7'b100_0000; // 0
		HEX2 <= 7'b000_0010; // 6
		end
		
		// 07 ~
		26'b00000000000000000001000000: begin
		HEX1 <= 7'b100_0000; // 0
		HEX2 <= 7'b111_1000; // 7
		end
		
		// 08 ~
		26'b00000000000000000010000000: begin
		HEX1 <= 7'b100_0000; // 0
		HEX2 <= 7'b000_0000; // 8
		end
		
		// 09 ~
		26'b00000000000000000100000000: begin
		HEX1 <= 7'b100_0000; // 0
		HEX2 <= 7'b001_1000; // 9
		end
		
		// 10 ~
		26'b00000000000000001000000000: begin
		HEX1 <= 7'b100_0000; // 0
		HEX2 <= 7'b000_1000; // A
		end
		
		// 11 ~
		26'b00000000000000010000000000: begin
		HEX1 <= 7'b100_0000; // 0
		HEX2 <= 7'b000_0011; // B
		end
		
		// 12 ~
		26'b00000000000000100000000000: begin
		HEX1 <= 7'b100_0000; // 0
		HEX2 <= 7'b100_0110; // C
		end
		
		// 13 ~
		26'b00000000000001000000000000: begin
		HEX1 <= 7'b100_0000; // 0
		HEX2 <= 7'b010_0001; // D
		end
		
		// 14 ~
		26'b00000000000010000000000000: begin
		HEX1 <= 7'b100_0000; // 0
		HEX2 <= 7'b000_0110; // E
		end
		
		// 15 ~
		26'b00000000000100000000000000: begin
		HEX1 <= 7'b100_0000; // 0
		HEX2 <= 7'b000_1110; // F
		end
		
		// 16 ~
		26'b00000000001000000000000000: begin
		HEX1 <= 7'b111_1001; // 1
		HEX2 <= 7'b100_0000; // 0
		end
		
		// 17 ~
		26'b00000000010000000000000000: begin
		HEX1 <= 7'b111_1001; // 1
		HEX2 <= 7'b111_1001; // 1
		end
		
		// 18 ~
		26'b00000000100000000000000000: begin
		HEX1 <= 7'b111_1001; // 1
		HEX2 <= 7'b010_0100; // 2
		end
		
		// 19 ~
		26'b00000001000000000000000000: begin
		HEX1 <= 7'b111_1001; // 1
		HEX2 <= 7'b011_0000; // 3
		end
		
		// 20 ~
		26'b00000010000000000000000000: begin
		HEX1 <= 7'b111_1001; // 1
		HEX2 <= 7'b001_1001; // 4
		end
		
		// 21 ~
		26'b00000100000000000000000000: begin
		HEX1 <= 7'b111_1001; // 1
		HEX2 <= 7'b001_0010; // 5
		end
		
		// 22 ~
		26'b00001000000000000000000000: begin
		HEX1 <= 7'b111_1001; // 1
		HEX2 <= 7'b000_0010; // 6
		end
		
		// 23 ~
		26'b00010000000000000000000000: begin
		HEX1 <= 7'b111_1001; // 1
		HEX2 <= 7'b111_1000; // 7
		end
		
		// 24 ~
		26'b00100000000000000000000000: begin
		HEX1 <= 7'b111_1001; // 1
		HEX2 <= 7'b000_0000; // 8
		end
		
		// 25 ~
		26'b01000000000000000000000000: begin
		HEX1 <= 7'b111_1001; // 1
		HEX2 <= 7'b001_1000; // 9
		end
		
		// 26 ~
		26'b10000000000000000000000000: begin
		HEX1 <= 7'b111_1001; // 1
		HEX2 <= 7'b000_1000; // A
		end
		
		//26'b01000000000000000000000000: HEX1 = 7'b100_0000 & HEX2 = 7'b010_0100;
		/*
		
		26'b10000000000000000000000000: begin
		HEX1 = 7'b111_1001;  HEX2 = 7'b010_0100;
		end
		
		//                 gfe_dcba
		4'b0000000000000000 : HEX = 7'b100_0000; // 0
		4'b0001 : HEX = 7'b111_1001; // 1
		4'b0010 : HEX = 7'b010_0100; // 2
		4'b0011 : HEX = 7'b011_0000; // 3
		4'b0100 : HEX = 7'b001_1001; // 4    
		4'b0101 : HEX = 7'b001_0010; // 5
		4'b0110 : HEX = 7'b000_0010; // 6
		4'b0111 : HEX = 7'b111_1000; // 7
		4'b1000 : HEX = 7'b000_0000; // 8
		4'b1001 : HEX = 7'b001_1000; // 9
		4'b1010 : HEX = 7'b000_1000; // A -> 10
		4'b1011 : HEX = 7'b000_0011; // B -> 11
		4'b1100 : HEX = 7'b100_0110; // C -> 12
		4'b1101 : HEX = 7'b010_0001; // D -> 13      
		4'b1110 : HEX = 7'b000_0110; // E -> 14
		4'b1111 : HEX = 7'b000_1110; // F -> 15
		
		default : HEX = 7'b000_0000; // Default Required
		*/
		default : begin 
		HEX1 <= 7'b000_0000; // Default Required
		HEX2 <= 7'b000_0000;
		end
		// Testing Vim commands
		endcase
	
endmodule

